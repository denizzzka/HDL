module tests;
    full_adder_test fa;
    alu_test a;
    nibble_counter_test nc;
    loopOverAllNibbles_test lan;
endmodule
