module tests;
    full_adder_test fa;
    loopOverAllNibbles_test lan;
endmodule
