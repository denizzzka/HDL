module tests;
    full_adder_test fa;
    alu_test a;
    loopOverAllNibbles_test lan;
    control_test c;
endmodule
